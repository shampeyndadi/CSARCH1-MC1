module MC1(F, A, B, C, D);
    hello
endmodule